module dff(d,clk,q,qbar);
input d,clk;
output  q ; 
output  qbar ;
 `include "dff_task.v"
always @(clk) begin
    dff_y(d,q,qbar);
end
endmodule